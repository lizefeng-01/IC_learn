typedef enum logic [1:0] {IDLE, S1, S2} state_t;

state_t state;
