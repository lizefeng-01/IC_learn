`include "uvm_macros.svh"
import uvm_pkg::*;


module top;
    initial begin
        run_test("my_test");
    end
endmodule




