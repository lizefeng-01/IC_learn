module tb_day5;

    bus_seq seq;

    initial begin
        seq = new();
        seq.run();
    end

endmodule
